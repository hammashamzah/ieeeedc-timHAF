library verilog;
use verilog.vl_types.all;
entity LUT_tb is
    port(
        theta           : out    vl_logic_vector(8 downto 0)
    );
end LUT_tb;
