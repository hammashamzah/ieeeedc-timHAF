module LUT(clock,code,theta);
    parameter n = 87;
    input         clock;
    input   [7:0] code;
    output  [7:0] theta;

    reg [7:0] theta;
    reg [7:0] code_in;

    always @(posedge clock)
        code_in <= code;

    always @(code_in)
    case(code_in)
        (8'd0): theta = 8'd90;
        (8'd1): theta = 8'd89;
        (8'd2): theta = 8'd89;
        (8'd3): theta = 8'd88;
        (8'd4): theta = 8'd87;
        (8'd5): theta = 8'd87;
        (8'd6): theta = 8'd86;
        (8'd7): theta = 8'd85;
        (8'd8): theta = 8'd85;
        (8'd9): theta = 8'd84;
        (8'd10): theta = 8'd83;
        (8'd11): theta = 8'd83;
        (8'd12): theta = 8'd82;
        (8'd13): theta = 8'd81;
        (8'd14): theta = 8'd81;
        (8'd15): theta = 8'd80;
        (8'd16): theta = 8'd79;
        (8'd17): theta = 8'd79;
        (8'd18): theta = 8'd78;
        (8'd19): theta = 8'd77;
        (8'd20): theta = 8'd77;
        (8'd21): theta = 8'd76;
        (8'd22): theta = 8'd75;
        (8'd23): theta = 8'd75;
        (8'd24): theta = 8'd74;
        (8'd25): theta = 8'd73;
        (8'd26): theta = 8'd73;
        (8'd27): theta = 8'd72;
        (8'd28): theta = 8'd71;
        (8'd29): theta = 8'd71;
        (8'd30): theta = 8'd70;
        (8'd31): theta = 8'd69;
        (8'd32): theta = 8'd68;
        (8'd33): theta = 8'd68;
        (8'd34): theta = 8'd67;
        (8'd35): theta = 8'd66;
        (8'd36): theta = 8'd66;
        (8'd37): theta = 8'd65;
        (8'd38): theta = 8'd64;
        (8'd39): theta = 8'd63;
        (8'd40): theta = 8'd63;
        (8'd41): theta = 8'd62;
        (8'd42): theta = 8'd61;
        (8'd43): theta = 8'd60;
        (8'd44): theta = 8'd60;
        (8'd45): theta = 8'd59;
        (8'd46): theta = 8'd58;
        (8'd47): theta = 8'd57;
        (8'd48): theta = 8'd56;
        (8'd49): theta = 8'd56;
        (8'd50): theta = 8'd55;
        (8'd51): theta = 8'd54;
        (8'd52): theta = 8'd53;
        (8'd53): theta = 8'd52;
        (8'd54): theta = 8'd52;
        (8'd55): theta = 8'd51;
        (8'd56): theta = 8'd50;
        (8'd57): theta = 8'd49;
        (8'd58): theta = 8'd48;
        (8'd59): theta = 8'd47;
        (8'd60): theta = 8'd46;
        (8'd61): theta = 8'd45;
        (8'd62): theta = 8'd45;
        (8'd63): theta = 8'd44;
        (8'd64): theta = 8'd43;
        (8'd65): theta = 8'd42;
        (8'd66): theta = 8'd41;
        (8'd67): theta = 8'd40;
        (8'd68): theta = 8'd39;
        (8'd69): theta = 8'd37;
        (8'd70): theta = 8'd36;
        (8'd71): theta = 8'd35;
        (8'd72): theta = 8'd34;
        (8'd73): theta = 8'd33;
        (8'd74): theta = 8'd32;
        (8'd75): theta = 8'd30;
        (8'd76): theta = 8'd29;
        (8'd77): theta = 8'd28;
        (8'd78): theta = 8'd26;
        (8'd79): theta = 8'd25;
        (8'd80): theta = 8'd23;
        (8'd81): theta = 8'd21;
        (8'd82): theta = 8'd19;
        (8'd83): theta = 8'd17;
        (8'd84): theta = 8'd15;
        (8'd85): theta = 8'd12;
        (8'd86): theta = 8'd9;
        default : theta = 8'd0;
    endcase
endmodule 