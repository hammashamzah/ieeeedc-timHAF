module LUT(clock,code,theta);
    parameter n = 87;
    input         clock;
    input   [6:0] code;
    output  [6:0] theta;

    reg [6:0] theta;
    reg [6:0] code_in;

    always @(posedge clock)
        code_in <= code;

    always @(code_in)
    case(code_in)
        (7'd0): theta = 7'd90;
        (7'd1): theta = 7'd89;
        (7'd2): theta = 7'd89;
        (7'd3): theta = 7'd88;
        (7'd4): theta = 7'd87;
        (7'd5): theta = 7'd87;
        (7'd6): theta = 7'd86;
        (7'd7): theta = 7'd85;
        (7'd8): theta = 7'd85;
        (7'd9): theta = 7'd84;
        (7'd10): theta = 7'd83;
        (7'd11): theta = 7'd83;
        (7'd12): theta = 7'd82;
        (7'd13): theta = 7'd81;
        (7'd14): theta = 7'd81;
        (7'd15): theta = 7'd80;
        (7'd16): theta = 7'd79;
        (7'd17): theta = 7'd79;
        (7'd18): theta = 7'd78;
        (7'd19): theta = 7'd77;
        (7'd20): theta = 7'd77;
        (7'd21): theta = 7'd76;
        (7'd22): theta = 7'd75;
        (7'd23): theta = 7'd75;
        (7'd24): theta = 7'd74;
        (7'd25): theta = 7'd73;
        (7'd26): theta = 7'd73;
        (7'd27): theta = 7'd72;
        (7'd28): theta = 7'd71;
        (7'd29): theta = 7'd71;
        (7'd30): theta = 7'd70;
        (7'd31): theta = 7'd69;
        (7'd32): theta = 7'd68;
        (7'd33): theta = 7'd68;
        (7'd34): theta = 7'd67;
        (7'd35): theta = 7'd66;
        (7'd36): theta = 7'd66;
        (7'd37): theta = 7'd65;
        (7'd38): theta = 7'd64;
        (7'd39): theta = 7'd63;
        (7'd40): theta = 7'd63;
        (7'd41): theta = 7'd62;
        (7'd42): theta = 7'd61;
        (7'd43): theta = 7'd60;
        (7'd44): theta = 7'd60;
        (7'd45): theta = 7'd59;
        (7'd46): theta = 7'd58;
        (7'd47): theta = 7'd57;
        (7'd48): theta = 7'd56;
        (7'd49): theta = 7'd56;
        (7'd50): theta = 7'd55;
        (7'd51): theta = 7'd54;
        (7'd52): theta = 7'd53;
        (7'd53): theta = 7'd52;
        (7'd54): theta = 7'd52;
        (7'd55): theta = 7'd51;
        (7'd56): theta = 7'd50;
        (7'd57): theta = 7'd49;
        (7'd58): theta = 7'd48;
        (7'd59): theta = 7'd47;
        (7'd60): theta = 7'd46;
        (7'd61): theta = 7'd45;
        (7'd62): theta = 7'd45;
        (7'd63): theta = 7'd44;
        (7'd64): theta = 7'd43;
        (7'd65): theta = 7'd42;
        (7'd66): theta = 7'd41;
        (7'd67): theta = 7'd40;
        (7'd68): theta = 7'd39;
        (7'd69): theta = 7'd37;
        (7'd70): theta = 7'd36;
        (7'd71): theta = 7'd35;
        (7'd72): theta = 7'd34;
        (7'd73): theta = 7'd33;
        (7'd74): theta = 7'd32;
        (7'd75): theta = 7'd30;
        (7'd76): theta = 7'd29;
        (7'd77): theta = 7'd28;
        (7'd78): theta = 7'd26;
        (7'd79): theta = 7'd25;
        (7'd80): theta = 7'd23;
        (7'd81): theta = 7'd21;
        (7'd82): theta = 7'd19;
        (7'd83): theta = 7'd17;
        (7'd84): theta = 7'd15;
        (7'd85): theta = 7'd12;
        (7'd86): theta = 7'd9;
        default : theta = 7'd0;
    endcase
endmodule 
